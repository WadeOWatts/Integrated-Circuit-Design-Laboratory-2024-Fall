# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : process_temp_1
#       Words            : 256
#       Bits             : 8
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2024/10/12 17:05:59
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO process_temp_1
CLASS BLOCK ;
FOREIGN process_temp_1 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 203.360 BY 215.600 ;
SYMMETRY x y r90 ;
SITE core_5040 ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 202.240 204.180 203.360 207.420 ;
  LAYER metal3 ;
  RECT 202.240 204.180 203.360 207.420 ;
  LAYER metal2 ;
  RECT 202.240 204.180 203.360 207.420 ;
  LAYER metal1 ;
  RECT 202.240 204.180 203.360 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 196.340 203.360 199.580 ;
  LAYER metal3 ;
  RECT 202.240 196.340 203.360 199.580 ;
  LAYER metal2 ;
  RECT 202.240 196.340 203.360 199.580 ;
  LAYER metal1 ;
  RECT 202.240 196.340 203.360 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 188.500 203.360 191.740 ;
  LAYER metal3 ;
  RECT 202.240 188.500 203.360 191.740 ;
  LAYER metal2 ;
  RECT 202.240 188.500 203.360 191.740 ;
  LAYER metal1 ;
  RECT 202.240 188.500 203.360 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 180.660 203.360 183.900 ;
  LAYER metal3 ;
  RECT 202.240 180.660 203.360 183.900 ;
  LAYER metal2 ;
  RECT 202.240 180.660 203.360 183.900 ;
  LAYER metal1 ;
  RECT 202.240 180.660 203.360 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 172.820 203.360 176.060 ;
  LAYER metal3 ;
  RECT 202.240 172.820 203.360 176.060 ;
  LAYER metal2 ;
  RECT 202.240 172.820 203.360 176.060 ;
  LAYER metal1 ;
  RECT 202.240 172.820 203.360 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 164.980 203.360 168.220 ;
  LAYER metal3 ;
  RECT 202.240 164.980 203.360 168.220 ;
  LAYER metal2 ;
  RECT 202.240 164.980 203.360 168.220 ;
  LAYER metal1 ;
  RECT 202.240 164.980 203.360 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 125.780 203.360 129.020 ;
  LAYER metal3 ;
  RECT 202.240 125.780 203.360 129.020 ;
  LAYER metal2 ;
  RECT 202.240 125.780 203.360 129.020 ;
  LAYER metal1 ;
  RECT 202.240 125.780 203.360 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 117.940 203.360 121.180 ;
  LAYER metal3 ;
  RECT 202.240 117.940 203.360 121.180 ;
  LAYER metal2 ;
  RECT 202.240 117.940 203.360 121.180 ;
  LAYER metal1 ;
  RECT 202.240 117.940 203.360 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 110.100 203.360 113.340 ;
  LAYER metal3 ;
  RECT 202.240 110.100 203.360 113.340 ;
  LAYER metal2 ;
  RECT 202.240 110.100 203.360 113.340 ;
  LAYER metal1 ;
  RECT 202.240 110.100 203.360 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 102.260 203.360 105.500 ;
  LAYER metal3 ;
  RECT 202.240 102.260 203.360 105.500 ;
  LAYER metal2 ;
  RECT 202.240 102.260 203.360 105.500 ;
  LAYER metal1 ;
  RECT 202.240 102.260 203.360 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 94.420 203.360 97.660 ;
  LAYER metal3 ;
  RECT 202.240 94.420 203.360 97.660 ;
  LAYER metal2 ;
  RECT 202.240 94.420 203.360 97.660 ;
  LAYER metal1 ;
  RECT 202.240 94.420 203.360 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 86.580 203.360 89.820 ;
  LAYER metal3 ;
  RECT 202.240 86.580 203.360 89.820 ;
  LAYER metal2 ;
  RECT 202.240 86.580 203.360 89.820 ;
  LAYER metal1 ;
  RECT 202.240 86.580 203.360 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 47.380 203.360 50.620 ;
  LAYER metal3 ;
  RECT 202.240 47.380 203.360 50.620 ;
  LAYER metal2 ;
  RECT 202.240 47.380 203.360 50.620 ;
  LAYER metal1 ;
  RECT 202.240 47.380 203.360 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 39.540 203.360 42.780 ;
  LAYER metal3 ;
  RECT 202.240 39.540 203.360 42.780 ;
  LAYER metal2 ;
  RECT 202.240 39.540 203.360 42.780 ;
  LAYER metal1 ;
  RECT 202.240 39.540 203.360 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 31.700 203.360 34.940 ;
  LAYER metal3 ;
  RECT 202.240 31.700 203.360 34.940 ;
  LAYER metal2 ;
  RECT 202.240 31.700 203.360 34.940 ;
  LAYER metal1 ;
  RECT 202.240 31.700 203.360 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 23.860 203.360 27.100 ;
  LAYER metal3 ;
  RECT 202.240 23.860 203.360 27.100 ;
  LAYER metal2 ;
  RECT 202.240 23.860 203.360 27.100 ;
  LAYER metal1 ;
  RECT 202.240 23.860 203.360 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 16.020 203.360 19.260 ;
  LAYER metal3 ;
  RECT 202.240 16.020 203.360 19.260 ;
  LAYER metal2 ;
  RECT 202.240 16.020 203.360 19.260 ;
  LAYER metal1 ;
  RECT 202.240 16.020 203.360 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 8.180 203.360 11.420 ;
  LAYER metal3 ;
  RECT 202.240 8.180 203.360 11.420 ;
  LAYER metal2 ;
  RECT 202.240 8.180 203.360 11.420 ;
  LAYER metal1 ;
  RECT 202.240 8.180 203.360 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 190.120 214.480 193.660 215.600 ;
  LAYER metal3 ;
  RECT 190.120 214.480 193.660 215.600 ;
  LAYER metal2 ;
  RECT 190.120 214.480 193.660 215.600 ;
  LAYER metal1 ;
  RECT 190.120 214.480 193.660 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 181.440 214.480 184.980 215.600 ;
  LAYER metal3 ;
  RECT 181.440 214.480 184.980 215.600 ;
  LAYER metal2 ;
  RECT 181.440 214.480 184.980 215.600 ;
  LAYER metal1 ;
  RECT 181.440 214.480 184.980 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 138.040 214.480 141.580 215.600 ;
  LAYER metal3 ;
  RECT 138.040 214.480 141.580 215.600 ;
  LAYER metal2 ;
  RECT 138.040 214.480 141.580 215.600 ;
  LAYER metal1 ;
  RECT 138.040 214.480 141.580 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 129.360 214.480 132.900 215.600 ;
  LAYER metal3 ;
  RECT 129.360 214.480 132.900 215.600 ;
  LAYER metal2 ;
  RECT 129.360 214.480 132.900 215.600 ;
  LAYER metal1 ;
  RECT 129.360 214.480 132.900 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 120.680 214.480 124.220 215.600 ;
  LAYER metal3 ;
  RECT 120.680 214.480 124.220 215.600 ;
  LAYER metal2 ;
  RECT 120.680 214.480 124.220 215.600 ;
  LAYER metal1 ;
  RECT 120.680 214.480 124.220 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 112.000 214.480 115.540 215.600 ;
  LAYER metal3 ;
  RECT 112.000 214.480 115.540 215.600 ;
  LAYER metal2 ;
  RECT 112.000 214.480 115.540 215.600 ;
  LAYER metal1 ;
  RECT 112.000 214.480 115.540 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 103.320 214.480 106.860 215.600 ;
  LAYER metal3 ;
  RECT 103.320 214.480 106.860 215.600 ;
  LAYER metal2 ;
  RECT 103.320 214.480 106.860 215.600 ;
  LAYER metal1 ;
  RECT 103.320 214.480 106.860 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 94.640 214.480 98.180 215.600 ;
  LAYER metal3 ;
  RECT 94.640 214.480 98.180 215.600 ;
  LAYER metal2 ;
  RECT 94.640 214.480 98.180 215.600 ;
  LAYER metal1 ;
  RECT 94.640 214.480 98.180 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 51.240 214.480 54.780 215.600 ;
  LAYER metal3 ;
  RECT 51.240 214.480 54.780 215.600 ;
  LAYER metal2 ;
  RECT 51.240 214.480 54.780 215.600 ;
  LAYER metal1 ;
  RECT 51.240 214.480 54.780 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 42.560 214.480 46.100 215.600 ;
  LAYER metal3 ;
  RECT 42.560 214.480 46.100 215.600 ;
  LAYER metal2 ;
  RECT 42.560 214.480 46.100 215.600 ;
  LAYER metal1 ;
  RECT 42.560 214.480 46.100 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 33.880 214.480 37.420 215.600 ;
  LAYER metal3 ;
  RECT 33.880 214.480 37.420 215.600 ;
  LAYER metal2 ;
  RECT 33.880 214.480 37.420 215.600 ;
  LAYER metal1 ;
  RECT 33.880 214.480 37.420 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.200 214.480 28.740 215.600 ;
  LAYER metal3 ;
  RECT 25.200 214.480 28.740 215.600 ;
  LAYER metal2 ;
  RECT 25.200 214.480 28.740 215.600 ;
  LAYER metal1 ;
  RECT 25.200 214.480 28.740 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 16.520 214.480 20.060 215.600 ;
  LAYER metal3 ;
  RECT 16.520 214.480 20.060 215.600 ;
  LAYER metal2 ;
  RECT 16.520 214.480 20.060 215.600 ;
  LAYER metal1 ;
  RECT 16.520 214.480 20.060 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.840 214.480 11.380 215.600 ;
  LAYER metal3 ;
  RECT 7.840 214.480 11.380 215.600 ;
  LAYER metal2 ;
  RECT 7.840 214.480 11.380 215.600 ;
  LAYER metal1 ;
  RECT 7.840 214.480 11.380 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 113.240 0.000 116.780 1.120 ;
  LAYER metal3 ;
  RECT 113.240 0.000 116.780 1.120 ;
  LAYER metal2 ;
  RECT 113.240 0.000 116.780 1.120 ;
  LAYER metal1 ;
  RECT 113.240 0.000 116.780 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 104.560 0.000 108.100 1.120 ;
  LAYER metal3 ;
  RECT 104.560 0.000 108.100 1.120 ;
  LAYER metal2 ;
  RECT 104.560 0.000 108.100 1.120 ;
  LAYER metal1 ;
  RECT 104.560 0.000 108.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 76.660 0.000 80.200 1.120 ;
  LAYER metal3 ;
  RECT 76.660 0.000 80.200 1.120 ;
  LAYER metal2 ;
  RECT 76.660 0.000 80.200 1.120 ;
  LAYER metal1 ;
  RECT 76.660 0.000 80.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 202.240 200.260 203.360 203.500 ;
  LAYER metal3 ;
  RECT 202.240 200.260 203.360 203.500 ;
  LAYER metal2 ;
  RECT 202.240 200.260 203.360 203.500 ;
  LAYER metal1 ;
  RECT 202.240 200.260 203.360 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 192.420 203.360 195.660 ;
  LAYER metal3 ;
  RECT 202.240 192.420 203.360 195.660 ;
  LAYER metal2 ;
  RECT 202.240 192.420 203.360 195.660 ;
  LAYER metal1 ;
  RECT 202.240 192.420 203.360 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 184.580 203.360 187.820 ;
  LAYER metal3 ;
  RECT 202.240 184.580 203.360 187.820 ;
  LAYER metal2 ;
  RECT 202.240 184.580 203.360 187.820 ;
  LAYER metal1 ;
  RECT 202.240 184.580 203.360 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 176.740 203.360 179.980 ;
  LAYER metal3 ;
  RECT 202.240 176.740 203.360 179.980 ;
  LAYER metal2 ;
  RECT 202.240 176.740 203.360 179.980 ;
  LAYER metal1 ;
  RECT 202.240 176.740 203.360 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 168.900 203.360 172.140 ;
  LAYER metal3 ;
  RECT 202.240 168.900 203.360 172.140 ;
  LAYER metal2 ;
  RECT 202.240 168.900 203.360 172.140 ;
  LAYER metal1 ;
  RECT 202.240 168.900 203.360 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 129.700 203.360 132.940 ;
  LAYER metal3 ;
  RECT 202.240 129.700 203.360 132.940 ;
  LAYER metal2 ;
  RECT 202.240 129.700 203.360 132.940 ;
  LAYER metal1 ;
  RECT 202.240 129.700 203.360 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 121.860 203.360 125.100 ;
  LAYER metal3 ;
  RECT 202.240 121.860 203.360 125.100 ;
  LAYER metal2 ;
  RECT 202.240 121.860 203.360 125.100 ;
  LAYER metal1 ;
  RECT 202.240 121.860 203.360 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 114.020 203.360 117.260 ;
  LAYER metal3 ;
  RECT 202.240 114.020 203.360 117.260 ;
  LAYER metal2 ;
  RECT 202.240 114.020 203.360 117.260 ;
  LAYER metal1 ;
  RECT 202.240 114.020 203.360 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 106.180 203.360 109.420 ;
  LAYER metal3 ;
  RECT 202.240 106.180 203.360 109.420 ;
  LAYER metal2 ;
  RECT 202.240 106.180 203.360 109.420 ;
  LAYER metal1 ;
  RECT 202.240 106.180 203.360 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 98.340 203.360 101.580 ;
  LAYER metal3 ;
  RECT 202.240 98.340 203.360 101.580 ;
  LAYER metal2 ;
  RECT 202.240 98.340 203.360 101.580 ;
  LAYER metal1 ;
  RECT 202.240 98.340 203.360 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 90.500 203.360 93.740 ;
  LAYER metal3 ;
  RECT 202.240 90.500 203.360 93.740 ;
  LAYER metal2 ;
  RECT 202.240 90.500 203.360 93.740 ;
  LAYER metal1 ;
  RECT 202.240 90.500 203.360 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 51.300 203.360 54.540 ;
  LAYER metal3 ;
  RECT 202.240 51.300 203.360 54.540 ;
  LAYER metal2 ;
  RECT 202.240 51.300 203.360 54.540 ;
  LAYER metal1 ;
  RECT 202.240 51.300 203.360 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 43.460 203.360 46.700 ;
  LAYER metal3 ;
  RECT 202.240 43.460 203.360 46.700 ;
  LAYER metal2 ;
  RECT 202.240 43.460 203.360 46.700 ;
  LAYER metal1 ;
  RECT 202.240 43.460 203.360 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 35.620 203.360 38.860 ;
  LAYER metal3 ;
  RECT 202.240 35.620 203.360 38.860 ;
  LAYER metal2 ;
  RECT 202.240 35.620 203.360 38.860 ;
  LAYER metal1 ;
  RECT 202.240 35.620 203.360 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 27.780 203.360 31.020 ;
  LAYER metal3 ;
  RECT 202.240 27.780 203.360 31.020 ;
  LAYER metal2 ;
  RECT 202.240 27.780 203.360 31.020 ;
  LAYER metal1 ;
  RECT 202.240 27.780 203.360 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 19.940 203.360 23.180 ;
  LAYER metal3 ;
  RECT 202.240 19.940 203.360 23.180 ;
  LAYER metal2 ;
  RECT 202.240 19.940 203.360 23.180 ;
  LAYER metal1 ;
  RECT 202.240 19.940 203.360 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 202.240 12.100 203.360 15.340 ;
  LAYER metal3 ;
  RECT 202.240 12.100 203.360 15.340 ;
  LAYER metal2 ;
  RECT 202.240 12.100 203.360 15.340 ;
  LAYER metal1 ;
  RECT 202.240 12.100 203.360 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 185.780 214.480 189.320 215.600 ;
  LAYER metal3 ;
  RECT 185.780 214.480 189.320 215.600 ;
  LAYER metal2 ;
  RECT 185.780 214.480 189.320 215.600 ;
  LAYER metal1 ;
  RECT 185.780 214.480 189.320 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 142.380 214.480 145.920 215.600 ;
  LAYER metal3 ;
  RECT 142.380 214.480 145.920 215.600 ;
  LAYER metal2 ;
  RECT 142.380 214.480 145.920 215.600 ;
  LAYER metal1 ;
  RECT 142.380 214.480 145.920 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 133.700 214.480 137.240 215.600 ;
  LAYER metal3 ;
  RECT 133.700 214.480 137.240 215.600 ;
  LAYER metal2 ;
  RECT 133.700 214.480 137.240 215.600 ;
  LAYER metal1 ;
  RECT 133.700 214.480 137.240 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 125.020 214.480 128.560 215.600 ;
  LAYER metal3 ;
  RECT 125.020 214.480 128.560 215.600 ;
  LAYER metal2 ;
  RECT 125.020 214.480 128.560 215.600 ;
  LAYER metal1 ;
  RECT 125.020 214.480 128.560 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 116.340 214.480 119.880 215.600 ;
  LAYER metal3 ;
  RECT 116.340 214.480 119.880 215.600 ;
  LAYER metal2 ;
  RECT 116.340 214.480 119.880 215.600 ;
  LAYER metal1 ;
  RECT 116.340 214.480 119.880 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 107.660 214.480 111.200 215.600 ;
  LAYER metal3 ;
  RECT 107.660 214.480 111.200 215.600 ;
  LAYER metal2 ;
  RECT 107.660 214.480 111.200 215.600 ;
  LAYER metal1 ;
  RECT 107.660 214.480 111.200 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 98.980 214.480 102.520 215.600 ;
  LAYER metal3 ;
  RECT 98.980 214.480 102.520 215.600 ;
  LAYER metal2 ;
  RECT 98.980 214.480 102.520 215.600 ;
  LAYER metal1 ;
  RECT 98.980 214.480 102.520 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 55.580 214.480 59.120 215.600 ;
  LAYER metal3 ;
  RECT 55.580 214.480 59.120 215.600 ;
  LAYER metal2 ;
  RECT 55.580 214.480 59.120 215.600 ;
  LAYER metal1 ;
  RECT 55.580 214.480 59.120 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 46.900 214.480 50.440 215.600 ;
  LAYER metal3 ;
  RECT 46.900 214.480 50.440 215.600 ;
  LAYER metal2 ;
  RECT 46.900 214.480 50.440 215.600 ;
  LAYER metal1 ;
  RECT 46.900 214.480 50.440 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 38.220 214.480 41.760 215.600 ;
  LAYER metal3 ;
  RECT 38.220 214.480 41.760 215.600 ;
  LAYER metal2 ;
  RECT 38.220 214.480 41.760 215.600 ;
  LAYER metal1 ;
  RECT 38.220 214.480 41.760 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 29.540 214.480 33.080 215.600 ;
  LAYER metal3 ;
  RECT 29.540 214.480 33.080 215.600 ;
  LAYER metal2 ;
  RECT 29.540 214.480 33.080 215.600 ;
  LAYER metal1 ;
  RECT 29.540 214.480 33.080 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 20.860 214.480 24.400 215.600 ;
  LAYER metal3 ;
  RECT 20.860 214.480 24.400 215.600 ;
  LAYER metal2 ;
  RECT 20.860 214.480 24.400 215.600 ;
  LAYER metal1 ;
  RECT 20.860 214.480 24.400 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.180 214.480 15.720 215.600 ;
  LAYER metal3 ;
  RECT 12.180 214.480 15.720 215.600 ;
  LAYER metal2 ;
  RECT 12.180 214.480 15.720 215.600 ;
  LAYER metal1 ;
  RECT 12.180 214.480 15.720 215.600 ;
 END
 PORT
  LAYER metal4 ;
  RECT 117.580 0.000 121.120 1.120 ;
  LAYER metal3 ;
  RECT 117.580 0.000 121.120 1.120 ;
  LAYER metal2 ;
  RECT 117.580 0.000 121.120 1.120 ;
  LAYER metal1 ;
  RECT 117.580 0.000 121.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 108.900 0.000 112.440 1.120 ;
  LAYER metal3 ;
  RECT 108.900 0.000 112.440 1.120 ;
  LAYER metal2 ;
  RECT 108.900 0.000 112.440 1.120 ;
  LAYER metal1 ;
  RECT 108.900 0.000 112.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 87.200 0.000 90.740 1.120 ;
  LAYER metal3 ;
  RECT 87.200 0.000 90.740 1.120 ;
  LAYER metal2 ;
  RECT 87.200 0.000 90.740 1.120 ;
  LAYER metal1 ;
  RECT 87.200 0.000 90.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 65.500 0.000 69.040 1.120 ;
  LAYER metal3 ;
  RECT 65.500 0.000 69.040 1.120 ;
  LAYER metal2 ;
  RECT 65.500 0.000 69.040 1.120 ;
  LAYER metal1 ;
  RECT 65.500 0.000 69.040 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal3 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal2 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal1 ;
  RECT 181.100 0.000 182.220 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal3 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal2 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal1 ;
  RECT 176.140 0.000 177.260 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal3 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal2 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal1 ;
  RECT 168.080 0.000 169.200 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 160.020 0.000 161.140 1.120 ;
  LAYER metal3 ;
  RECT 160.020 0.000 161.140 1.120 ;
  LAYER metal2 ;
  RECT 160.020 0.000 161.140 1.120 ;
  LAYER metal1 ;
  RECT 160.020 0.000 161.140 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 151.340 0.000 152.460 1.120 ;
  LAYER metal3 ;
  RECT 151.340 0.000 152.460 1.120 ;
  LAYER metal2 ;
  RECT 151.340 0.000 152.460 1.120 ;
  LAYER metal1 ;
  RECT 151.340 0.000 152.460 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER metal3 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER metal2 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER metal1 ;
  RECT 138.320 0.000 139.440 1.120 ;
 END
END DI4
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 132.120 0.000 133.240 1.120 ;
  LAYER metal3 ;
  RECT 132.120 0.000 133.240 1.120 ;
  LAYER metal2 ;
  RECT 132.120 0.000 133.240 1.120 ;
  LAYER metal1 ;
  RECT 132.120 0.000 133.240 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 130.260 0.000 131.380 1.120 ;
  LAYER metal3 ;
  RECT 130.260 0.000 131.380 1.120 ;
  LAYER metal2 ;
  RECT 130.260 0.000 131.380 1.120 ;
  LAYER metal1 ;
  RECT 130.260 0.000 131.380 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER metal4 ;
  RECT 125.920 0.000 127.040 1.120 ;
  LAYER metal3 ;
  RECT 125.920 0.000 127.040 1.120 ;
  LAYER metal2 ;
  RECT 125.920 0.000 127.040 1.120 ;
  LAYER metal1 ;
  RECT 125.920 0.000 127.040 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER metal4 ;
  RECT 124.060 0.000 125.180 1.120 ;
  LAYER metal3 ;
  RECT 124.060 0.000 125.180 1.120 ;
  LAYER metal2 ;
  RECT 124.060 0.000 125.180 1.120 ;
  LAYER metal1 ;
  RECT 124.060 0.000 125.180 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 102.360 0.000 103.480 1.120 ;
  LAYER metal3 ;
  RECT 102.360 0.000 103.480 1.120 ;
  LAYER metal2 ;
  RECT 102.360 0.000 103.480 1.120 ;
  LAYER metal1 ;
  RECT 102.360 0.000 103.480 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER metal4 ;
  RECT 99.260 0.000 100.380 1.120 ;
  LAYER metal3 ;
  RECT 99.260 0.000 100.380 1.120 ;
  LAYER metal2 ;
  RECT 99.260 0.000 100.380 1.120 ;
  LAYER metal1 ;
  RECT 99.260 0.000 100.380 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 96.780 0.000 97.900 1.120 ;
  LAYER metal3 ;
  RECT 96.780 0.000 97.900 1.120 ;
  LAYER metal2 ;
  RECT 96.780 0.000 97.900 1.120 ;
  LAYER metal1 ;
  RECT 96.780 0.000 97.900 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 92.440 0.000 93.560 1.120 ;
  LAYER metal3 ;
  RECT 92.440 0.000 93.560 1.120 ;
  LAYER metal2 ;
  RECT 92.440 0.000 93.560 1.120 ;
  LAYER metal1 ;
  RECT 92.440 0.000 93.560 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 85.000 0.000 86.120 1.120 ;
  LAYER metal3 ;
  RECT 85.000 0.000 86.120 1.120 ;
  LAYER metal2 ;
  RECT 85.000 0.000 86.120 1.120 ;
  LAYER metal1 ;
  RECT 85.000 0.000 86.120 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 81.900 0.000 83.020 1.120 ;
  LAYER metal3 ;
  RECT 81.900 0.000 83.020 1.120 ;
  LAYER metal2 ;
  RECT 81.900 0.000 83.020 1.120 ;
  LAYER metal1 ;
  RECT 81.900 0.000 83.020 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 74.460 0.000 75.580 1.120 ;
  LAYER metal3 ;
  RECT 74.460 0.000 75.580 1.120 ;
  LAYER metal2 ;
  RECT 74.460 0.000 75.580 1.120 ;
  LAYER metal1 ;
  RECT 74.460 0.000 75.580 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 71.360 0.000 72.480 1.120 ;
  LAYER metal3 ;
  RECT 71.360 0.000 72.480 1.120 ;
  LAYER metal2 ;
  RECT 71.360 0.000 72.480 1.120 ;
  LAYER metal1 ;
  RECT 71.360 0.000 72.480 1.120 ;
 END
END A7
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 203.360 215.600 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 203.360 215.600 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 203.360 215.600 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 203.360 215.600 ;
  LAYER via ;
  RECT 0.000 0.140 203.360 215.600 ;
  LAYER via2 ;
  RECT 0.000 0.140 203.360 215.600 ;
  LAYER via3 ;
  RECT 0.000 0.140 203.360 215.600 ;
END
END process_temp_1
END LIBRARY



